-- disenyo_qsys_tb.vhd

-- Generated using ACDS version 19.1 670

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity disenyo_qsys_tb is
end entity disenyo_qsys_tb;

architecture rtl of disenyo_qsys_tb is
	component disenyo_qsys is
		port (
			clk_clk          : in    std_logic                     := 'X';             -- clk
			reset_reset_n    : in    std_logic                     := 'X';             -- reset_n
			sdram_clk_clk    : out   std_logic;                                        -- clk
			sdram_wire_addr  : out   std_logic_vector(12 downto 0);                    -- addr
			sdram_wire_ba    : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_wire_cas_n : out   std_logic;                                        -- cas_n
			sdram_wire_cke   : out   std_logic;                                        -- cke
			sdram_wire_cs_n  : out   std_logic;                                        -- cs_n
			sdram_wire_dq    : inout std_logic_vector(31 downto 0) := (others => 'X'); -- dq
			sdram_wire_dqm   : out   std_logic_vector(3 downto 0);                     -- dqm
			sdram_wire_ras_n : out   std_logic;                                        -- ras_n
			sdram_wire_we_n  : out   std_logic                                         -- we_n
		);
	end component disenyo_qsys;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_sdram_partner_module is
		port (
			clk      : in    std_logic                     := 'X';             -- clk
			zs_dq    : inout std_logic_vector(31 downto 0) := (others => 'X'); -- dq
			zs_addr  : in    std_logic_vector(12 downto 0) := (others => 'X'); -- addr
			zs_ba    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- ba
			zs_cas_n : in    std_logic                     := 'X';             -- cas_n
			zs_cke   : in    std_logic                     := 'X';             -- cke
			zs_cs_n  : in    std_logic                     := 'X';             -- cs_n
			zs_dqm   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- dqm
			zs_ras_n : in    std_logic                     := 'X';             -- ras_n
			zs_we_n  : in    std_logic                     := 'X'              -- we_n
		);
	end component altera_sdram_partner_module;

	signal disenyo_qsys_inst_clk_bfm_clk_clk                 : std_logic;                     -- disenyo_qsys_inst_clk_bfm:clk -> [disenyo_qsys_inst:clk_clk, disenyo_qsys_inst_reset_bfm:clk]
	signal new_sdram_controller_0_my_partner_clk_bfm_clk_clk : std_logic;                     -- new_sdram_controller_0_my_partner_clk_bfm:clk -> new_sdram_controller_0_my_partner:clk
	signal disenyo_qsys_inst_sdram_wire_cs_n                 : std_logic;                     -- disenyo_qsys_inst:sdram_wire_cs_n -> new_sdram_controller_0_my_partner:zs_cs_n
	signal disenyo_qsys_inst_sdram_wire_dqm                  : std_logic_vector(3 downto 0);  -- disenyo_qsys_inst:sdram_wire_dqm -> new_sdram_controller_0_my_partner:zs_dqm
	signal disenyo_qsys_inst_sdram_wire_cas_n                : std_logic;                     -- disenyo_qsys_inst:sdram_wire_cas_n -> new_sdram_controller_0_my_partner:zs_cas_n
	signal disenyo_qsys_inst_sdram_wire_ras_n                : std_logic;                     -- disenyo_qsys_inst:sdram_wire_ras_n -> new_sdram_controller_0_my_partner:zs_ras_n
	signal disenyo_qsys_inst_sdram_wire_we_n                 : std_logic;                     -- disenyo_qsys_inst:sdram_wire_we_n -> new_sdram_controller_0_my_partner:zs_we_n
	signal disenyo_qsys_inst_sdram_wire_addr                 : std_logic_vector(12 downto 0); -- disenyo_qsys_inst:sdram_wire_addr -> new_sdram_controller_0_my_partner:zs_addr
	signal disenyo_qsys_inst_sdram_wire_cke                  : std_logic;                     -- disenyo_qsys_inst:sdram_wire_cke -> new_sdram_controller_0_my_partner:zs_cke
	signal disenyo_qsys_inst_sdram_wire_dq                   : std_logic_vector(31 downto 0); -- [] -> [disenyo_qsys_inst:sdram_wire_dq, new_sdram_controller_0_my_partner:zs_dq]
	signal disenyo_qsys_inst_sdram_wire_ba                   : std_logic_vector(1 downto 0);  -- disenyo_qsys_inst:sdram_wire_ba -> new_sdram_controller_0_my_partner:zs_ba
	signal disenyo_qsys_inst_reset_bfm_reset_reset           : std_logic;                     -- disenyo_qsys_inst_reset_bfm:reset -> disenyo_qsys_inst:reset_reset_n

begin

	disenyo_qsys_inst : component disenyo_qsys
		port map (
			clk_clk          => disenyo_qsys_inst_clk_bfm_clk_clk,       --        clk.clk
			reset_reset_n    => disenyo_qsys_inst_reset_bfm_reset_reset, --      reset.reset_n
			sdram_clk_clk    => open,                                    --  sdram_clk.clk
			sdram_wire_addr  => disenyo_qsys_inst_sdram_wire_addr,       -- sdram_wire.addr
			sdram_wire_ba    => disenyo_qsys_inst_sdram_wire_ba,         --           .ba
			sdram_wire_cas_n => disenyo_qsys_inst_sdram_wire_cas_n,      --           .cas_n
			sdram_wire_cke   => disenyo_qsys_inst_sdram_wire_cke,        --           .cke
			sdram_wire_cs_n  => disenyo_qsys_inst_sdram_wire_cs_n,       --           .cs_n
			sdram_wire_dq    => disenyo_qsys_inst_sdram_wire_dq,         --           .dq
			sdram_wire_dqm   => disenyo_qsys_inst_sdram_wire_dqm,        --           .dqm
			sdram_wire_ras_n => disenyo_qsys_inst_sdram_wire_ras_n,      --           .ras_n
			sdram_wire_we_n  => disenyo_qsys_inst_sdram_wire_we_n        --           .we_n
		);

	disenyo_qsys_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => disenyo_qsys_inst_clk_bfm_clk_clk  -- clk.clk
		);

	disenyo_qsys_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => disenyo_qsys_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => disenyo_qsys_inst_clk_bfm_clk_clk        --   clk.clk
		);

	new_sdram_controller_0_my_partner : component altera_sdram_partner_module
		port map (
			clk      => new_sdram_controller_0_my_partner_clk_bfm_clk_clk, --     clk.clk
			zs_dq    => disenyo_qsys_inst_sdram_wire_dq,                   -- conduit.dq
			zs_addr  => disenyo_qsys_inst_sdram_wire_addr,                 --        .addr
			zs_ba    => disenyo_qsys_inst_sdram_wire_ba,                   --        .ba
			zs_cas_n => disenyo_qsys_inst_sdram_wire_cas_n,                --        .cas_n
			zs_cke   => disenyo_qsys_inst_sdram_wire_cke,                  --        .cke
			zs_cs_n  => disenyo_qsys_inst_sdram_wire_cs_n,                 --        .cs_n
			zs_dqm   => disenyo_qsys_inst_sdram_wire_dqm,                  --        .dqm
			zs_ras_n => disenyo_qsys_inst_sdram_wire_ras_n,                --        .ras_n
			zs_we_n  => disenyo_qsys_inst_sdram_wire_we_n                  --        .we_n
		);

	new_sdram_controller_0_my_partner_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => new_sdram_controller_0_my_partner_clk_bfm_clk_clk  -- clk.clk
		);

end architecture rtl; -- of disenyo_qsys_tb
