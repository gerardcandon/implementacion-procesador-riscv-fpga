-- disenyo_qsys.vhd

-- Generated using ACDS version 19.1 670

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity disenyo_qsys is
	port (
		clk_clk          : in    std_logic                     := '0';             --        clk.clk
		ps2_CLK          : inout std_logic                     := '0';             --        ps2.CLK
		ps2_DAT          : inout std_logic                     := '0';             --           .DAT
		reset_reset_n    : in    std_logic                     := '0';             --      reset.reset_n
		sdram_clk_clk    : out   std_logic;                                        --  sdram_clk.clk
		sdram_wire_addr  : out   std_logic_vector(12 downto 0);                    -- sdram_wire.addr
		sdram_wire_ba    : out   std_logic_vector(1 downto 0);                     --           .ba
		sdram_wire_cas_n : out   std_logic;                                        --           .cas_n
		sdram_wire_cke   : out   std_logic;                                        --           .cke
		sdram_wire_cs_n  : out   std_logic;                                        --           .cs_n
		sdram_wire_dq    : inout std_logic_vector(31 downto 0) := (others => '0'); --           .dq
		sdram_wire_dqm   : out   std_logic_vector(3 downto 0);                     --           .dqm
		sdram_wire_ras_n : out   std_logic;                                        --           .ras_n
		sdram_wire_we_n  : out   std_logic;                                        --           .we_n
		sram_DQ          : inout std_logic_vector(15 downto 0) := (others => '0'); --       sram.DQ
		sram_ADDR        : out   std_logic_vector(19 downto 0);                    --           .ADDR
		sram_LB_N        : out   std_logic;                                        --           .LB_N
		sram_UB_N        : out   std_logic;                                        --           .UB_N
		sram_CE_N        : out   std_logic;                                        --           .CE_N
		sram_OE_N        : out   std_logic;                                        --           .OE_N
		sram_WE_N        : out   std_logic;                                        --           .WE_N
		start_bit        : in    std_logic                     := '0';             --      start.bit
		vga_CLK          : out   std_logic;                                        --        vga.CLK
		vga_HS           : out   std_logic;                                        --           .HS
		vga_VS           : out   std_logic;                                        --           .VS
		vga_BLANK        : out   std_logic;                                        --           .BLANK
		vga_SYNC         : out   std_logic;                                        --           .SYNC
		vga_R            : out   std_logic_vector(7 downto 0);                     --           .R
		vga_G            : out   std_logic_vector(7 downto 0);                     --           .G
		vga_B            : out   std_logic_vector(7 downto 0)                      --           .B
	);
end entity disenyo_qsys;

architecture rtl of disenyo_qsys is
	component ensamblado_procesador is
		port (
			reset         : in  std_logic                     := 'X';             -- reset
			address       : out std_logic_vector(31 downto 0);                    -- address
			writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			read          : out std_logic;                                        -- read
			write         : out std_logic;                                        -- write
			byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			reloj         : in  std_logic                     := 'X';             -- clk
			irq           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- irq
			start         : in  std_logic                     := 'X'              -- bit
		);
	end component ensamblado_procesador;

	component disenyo_qsys_master_0 is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component disenyo_qsys_master_0;

	component mm_reloj is
		port (
			read          : in  std_logic                     := 'X';             -- read
			write         : in  std_logic                     := 'X';             -- write
			address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			waitrequest   : out std_logic;                                        -- waitrequest
			readdatavalid : out std_logic;                                        -- readdatavalid
			Pcero         : in  std_logic                     := 'X';             -- reset
			reloj         : in  std_logic                     := 'X';             -- clk
			int_clk       : out std_logic                                         -- irq
		);
	end component mm_reloj;

	component disenyo_qsys_new_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component disenyo_qsys_new_sdram_controller_0;

	component disenyo_qsys_ps2_0 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic                     := 'X';             -- address
			chipselect  : in    std_logic                     := 'X';             -- chipselect
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			irq         : out   std_logic;                                        -- irq
			PS2_CLK     : inout std_logic                     := 'X';             -- export
			PS2_DAT     : inout std_logic                     := 'X'              -- export
		);
	end component disenyo_qsys_ps2_0;

	component disenyo_qsys_sram_0 is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component disenyo_qsys_sram_0;

	component disenyo_qsys_sys_sdram_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component disenyo_qsys_sys_sdram_pll_0;

	component disenyo_qsys_video_dma_controller_0 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_data          : out std_logic_vector(29 downto 0);                    -- data
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic                                         -- valid
		);
	end component disenyo_qsys_video_dma_controller_0;

	component disenyo_qsys_video_dual_clock_buffer_0 is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component disenyo_qsys_video_dual_clock_buffer_0;

	component disenyo_qsys_video_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			vga_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component disenyo_qsys_video_pll_0;

	component disenyo_qsys_video_vga_controller_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(7 downto 0);                     -- export
			VGA_G         : out std_logic_vector(7 downto 0);                     -- export
			VGA_B         : out std_logic_vector(7 downto 0)                      -- export
		);
	end component disenyo_qsys_video_vga_controller_0;

	component disenyo_qsys_mm_interconnect_0 is
		port (
			sys_sdram_pll_0_sys_clk_clk                                : in  std_logic                     := 'X';             -- clk
			master_0_clk_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			new_sdram_controller_0_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			video_dma_controller_0_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			ensamblado_procesador_0_avalon_master_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			ensamblado_procesador_0_avalon_master_waitrequest          : out std_logic;                                        -- waitrequest
			ensamblado_procesador_0_avalon_master_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ensamblado_procesador_0_avalon_master_read                 : in  std_logic                     := 'X';             -- read
			ensamblado_procesador_0_avalon_master_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			ensamblado_procesador_0_avalon_master_readdatavalid        : out std_logic;                                        -- readdatavalid
			ensamblado_procesador_0_avalon_master_write                : in  std_logic                     := 'X';             -- write
			ensamblado_procesador_0_avalon_master_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			master_0_master_address                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			master_0_master_waitrequest                                : out std_logic;                                        -- waitrequest
			master_0_master_byteenable                                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			master_0_master_read                                       : in  std_logic                     := 'X';             -- read
			master_0_master_readdata                                   : out std_logic_vector(31 downto 0);                    -- readdata
			master_0_master_readdatavalid                              : out std_logic;                                        -- readdatavalid
			master_0_master_write                                      : in  std_logic                     := 'X';             -- write
			master_0_master_writedata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			video_dma_controller_0_avalon_dma_master_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			video_dma_controller_0_avalon_dma_master_waitrequest       : out std_logic;                                        -- waitrequest
			video_dma_controller_0_avalon_dma_master_read              : in  std_logic                     := 'X';             -- read
			video_dma_controller_0_avalon_dma_master_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			video_dma_controller_0_avalon_dma_master_readdatavalid     : out std_logic;                                        -- readdatavalid
			video_dma_controller_0_avalon_dma_master_lock              : in  std_logic                     := 'X';             -- lock
			mm_reloj_0_avalon_slave_0_address                          : out std_logic_vector(3 downto 0);                     -- address
			mm_reloj_0_avalon_slave_0_write                            : out std_logic;                                        -- write
			mm_reloj_0_avalon_slave_0_read                             : out std_logic;                                        -- read
			mm_reloj_0_avalon_slave_0_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mm_reloj_0_avalon_slave_0_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			mm_reloj_0_avalon_slave_0_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			mm_reloj_0_avalon_slave_0_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			mm_reloj_0_avalon_slave_0_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			new_sdram_controller_0_s1_address                          : out std_logic_vector(24 downto 0);                    -- address
			new_sdram_controller_0_s1_write                            : out std_logic;                                        -- write
			new_sdram_controller_0_s1_read                             : out std_logic;                                        -- read
			new_sdram_controller_0_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			new_sdram_controller_0_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			new_sdram_controller_0_s1_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			new_sdram_controller_0_s1_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			new_sdram_controller_0_s1_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			new_sdram_controller_0_s1_chipselect                       : out std_logic;                                        -- chipselect
			ps2_0_avalon_ps2_slave_address                             : out std_logic_vector(0 downto 0);                     -- address
			ps2_0_avalon_ps2_slave_write                               : out std_logic;                                        -- write
			ps2_0_avalon_ps2_slave_read                                : out std_logic;                                        -- read
			ps2_0_avalon_ps2_slave_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ps2_0_avalon_ps2_slave_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			ps2_0_avalon_ps2_slave_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			ps2_0_avalon_ps2_slave_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			ps2_0_avalon_ps2_slave_chipselect                          : out std_logic;                                        -- chipselect
			sram_0_avalon_sram_slave_address                           : out std_logic_vector(19 downto 0);                    -- address
			sram_0_avalon_sram_slave_write                             : out std_logic;                                        -- write
			sram_0_avalon_sram_slave_read                              : out std_logic;                                        -- read
			sram_0_avalon_sram_slave_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sram_0_avalon_sram_slave_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			sram_0_avalon_sram_slave_byteenable                        : out std_logic_vector(1 downto 0);                     -- byteenable
			sram_0_avalon_sram_slave_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			video_dma_controller_0_avalon_dma_control_slave_address    : out std_logic_vector(1 downto 0);                     -- address
			video_dma_controller_0_avalon_dma_control_slave_write      : out std_logic;                                        -- write
			video_dma_controller_0_avalon_dma_control_slave_read       : out std_logic;                                        -- read
			video_dma_controller_0_avalon_dma_control_slave_readdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			video_dma_controller_0_avalon_dma_control_slave_writedata  : out std_logic_vector(31 downto 0);                    -- writedata
			video_dma_controller_0_avalon_dma_control_slave_byteenable : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component disenyo_qsys_mm_interconnect_0;

	component disenyo_qsys_irq_mapper is
		port (
			clk           : in  std_logic                    := 'X'; -- clk
			reset         : in  std_logic                    := 'X'; -- reset
			receiver0_irq : in  std_logic                    := 'X'; -- irq
			receiver1_irq : in  std_logic                    := 'X'; -- irq
			sender_irq    : out std_logic_vector(1 downto 0)         -- irq
		);
	end component disenyo_qsys_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_valid                      : std_logic;                     -- video_dual_clock_buffer_0:stream_out_valid -> video_vga_controller_0:valid
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_data                       : std_logic_vector(29 downto 0); -- video_dual_clock_buffer_0:stream_out_data -> video_vga_controller_0:data
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_ready                      : std_logic;                     -- video_vga_controller_0:ready -> video_dual_clock_buffer_0:stream_out_ready
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket              : std_logic;                     -- video_dual_clock_buffer_0:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket                : std_logic;                     -- video_dual_clock_buffer_0:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	signal video_dma_controller_0_avalon_pixel_source_valid                             : std_logic;                     -- video_dma_controller_0:stream_valid -> video_dual_clock_buffer_0:stream_in_valid
	signal video_dma_controller_0_avalon_pixel_source_data                              : std_logic_vector(29 downto 0); -- video_dma_controller_0:stream_data -> video_dual_clock_buffer_0:stream_in_data
	signal video_dma_controller_0_avalon_pixel_source_ready                             : std_logic;                     -- video_dual_clock_buffer_0:stream_in_ready -> video_dma_controller_0:stream_ready
	signal video_dma_controller_0_avalon_pixel_source_startofpacket                     : std_logic;                     -- video_dma_controller_0:stream_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	signal video_dma_controller_0_avalon_pixel_source_endofpacket                       : std_logic;                     -- video_dma_controller_0:stream_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	signal sys_sdram_pll_0_sys_clk_clk                                                  : std_logic;                     -- sys_sdram_pll_0:sys_clk_clk -> [ensamblado_procesador_0:reloj, irq_mapper:clk, master_0:clk_clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, mm_reloj_0:reloj, new_sdram_controller_0:clk, ps2_0:clk, rst_controller:clk, rst_controller_001:clk, sram_0:clk, video_dma_controller_0:clk, video_dual_clock_buffer_0:clk_stream_in, video_pll_0:ref_clk_clk]
	signal video_pll_0_vga_clk_clk                                                      : std_logic;                     -- video_pll_0:vga_clk_clk -> [rst_controller_003:clk, video_dual_clock_buffer_0:clk_stream_out, video_vga_controller_0:clk]
	signal video_dma_controller_0_avalon_dma_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:video_dma_controller_0_avalon_dma_master_waitrequest -> video_dma_controller_0:master_waitrequest
	signal video_dma_controller_0_avalon_dma_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdata -> video_dma_controller_0:master_readdata
	signal video_dma_controller_0_avalon_dma_master_address                             : std_logic_vector(31 downto 0); -- video_dma_controller_0:master_address -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_address
	signal video_dma_controller_0_avalon_dma_master_read                                : std_logic;                     -- video_dma_controller_0:master_read -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_read
	signal video_dma_controller_0_avalon_dma_master_readdatavalid                       : std_logic;                     -- mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdatavalid -> video_dma_controller_0:master_readdatavalid
	signal video_dma_controller_0_avalon_dma_master_lock                                : std_logic;                     -- video_dma_controller_0:master_arbiterlock -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_lock
	signal ensamblado_procesador_0_avalon_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:ensamblado_procesador_0_avalon_master_readdata -> ensamblado_procesador_0:readdata
	signal ensamblado_procesador_0_avalon_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:ensamblado_procesador_0_avalon_master_waitrequest -> ensamblado_procesador_0:waitrequest
	signal ensamblado_procesador_0_avalon_master_address                                : std_logic_vector(31 downto 0); -- ensamblado_procesador_0:address -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_address
	signal ensamblado_procesador_0_avalon_master_read                                   : std_logic;                     -- ensamblado_procesador_0:read -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_read
	signal ensamblado_procesador_0_avalon_master_byteenable                             : std_logic_vector(3 downto 0);  -- ensamblado_procesador_0:byteenable -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_byteenable
	signal ensamblado_procesador_0_avalon_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:ensamblado_procesador_0_avalon_master_readdatavalid -> ensamblado_procesador_0:readdatavalid
	signal ensamblado_procesador_0_avalon_master_writedata                              : std_logic_vector(31 downto 0); -- ensamblado_procesador_0:writedata -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_writedata
	signal ensamblado_procesador_0_avalon_master_write                                  : std_logic;                     -- ensamblado_procesador_0:write -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_write
	signal master_0_master_readdata                                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	signal master_0_master_waitrequest                                                  : std_logic;                     -- mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	signal master_0_master_address                                                      : std_logic_vector(31 downto 0); -- master_0:master_address -> mm_interconnect_0:master_0_master_address
	signal master_0_master_read                                                         : std_logic;                     -- master_0:master_read -> mm_interconnect_0:master_0_master_read
	signal master_0_master_byteenable                                                   : std_logic_vector(3 downto 0);  -- master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	signal master_0_master_readdatavalid                                                : std_logic;                     -- mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	signal master_0_master_write                                                        : std_logic;                     -- master_0:master_write -> mm_interconnect_0:master_0_master_write
	signal master_0_master_writedata                                                    : std_logic_vector(31 downto 0); -- master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	signal mm_interconnect_0_sram_0_avalon_sram_slave_readdata                          : std_logic_vector(15 downto 0); -- sram_0:readdata -> mm_interconnect_0:sram_0_avalon_sram_slave_readdata
	signal mm_interconnect_0_sram_0_avalon_sram_slave_address                           : std_logic_vector(19 downto 0); -- mm_interconnect_0:sram_0_avalon_sram_slave_address -> sram_0:address
	signal mm_interconnect_0_sram_0_avalon_sram_slave_read                              : std_logic;                     -- mm_interconnect_0:sram_0_avalon_sram_slave_read -> sram_0:read
	signal mm_interconnect_0_sram_0_avalon_sram_slave_byteenable                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sram_0_avalon_sram_slave_byteenable -> sram_0:byteenable
	signal mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid                     : std_logic;                     -- sram_0:readdatavalid -> mm_interconnect_0:sram_0_avalon_sram_slave_readdatavalid
	signal mm_interconnect_0_sram_0_avalon_sram_slave_write                             : std_logic;                     -- mm_interconnect_0:sram_0_avalon_sram_slave_write -> sram_0:write
	signal mm_interconnect_0_sram_0_avalon_sram_slave_writedata                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:sram_0_avalon_sram_slave_writedata -> sram_0:writedata
	signal mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_readdata   : std_logic_vector(31 downto 0); -- video_dma_controller_0:slave_readdata -> mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_readdata
	signal mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_address -> video_dma_controller_0:slave_address
	signal mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_read       : std_logic;                     -- mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_read -> video_dma_controller_0:slave_read
	signal mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_byteenable -> video_dma_controller_0:slave_byteenable
	signal mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_write      : std_logic;                     -- mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_write -> video_dma_controller_0:slave_write
	signal mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_writedata -> video_dma_controller_0:slave_writedata
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_chipselect                          : std_logic;                     -- mm_interconnect_0:ps2_0_avalon_ps2_slave_chipselect -> ps2_0:chipselect
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_readdata                            : std_logic_vector(31 downto 0); -- ps2_0:readdata -> mm_interconnect_0:ps2_0_avalon_ps2_slave_readdata
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_waitrequest                         : std_logic;                     -- ps2_0:waitrequest -> mm_interconnect_0:ps2_0_avalon_ps2_slave_waitrequest
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_address                             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ps2_0_avalon_ps2_slave_address -> ps2_0:address
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_read                                : std_logic;                     -- mm_interconnect_0:ps2_0_avalon_ps2_slave_read -> ps2_0:read
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ps2_0_avalon_ps2_slave_byteenable -> ps2_0:byteenable
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_write                               : std_logic;                     -- mm_interconnect_0:ps2_0_avalon_ps2_slave_write -> ps2_0:write
	signal mm_interconnect_0_ps2_0_avalon_ps2_slave_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:ps2_0_avalon_ps2_slave_writedata -> ps2_0:writedata
	signal mm_interconnect_0_mm_reloj_0_avalon_slave_0_readdata                         : std_logic_vector(31 downto 0); -- mm_reloj_0:readdata -> mm_interconnect_0:mm_reloj_0_avalon_slave_0_readdata
	signal mm_interconnect_0_mm_reloj_0_avalon_slave_0_waitrequest                      : std_logic;                     -- mm_reloj_0:waitrequest -> mm_interconnect_0:mm_reloj_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_mm_reloj_0_avalon_slave_0_address                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:mm_reloj_0_avalon_slave_0_address -> mm_reloj_0:address
	signal mm_interconnect_0_mm_reloj_0_avalon_slave_0_read                             : std_logic;                     -- mm_interconnect_0:mm_reloj_0_avalon_slave_0_read -> mm_reloj_0:read
	signal mm_interconnect_0_mm_reloj_0_avalon_slave_0_byteenable                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:mm_reloj_0_avalon_slave_0_byteenable -> mm_reloj_0:byteenable
	signal mm_interconnect_0_mm_reloj_0_avalon_slave_0_readdatavalid                    : std_logic;                     -- mm_reloj_0:readdatavalid -> mm_interconnect_0:mm_reloj_0_avalon_slave_0_readdatavalid
	signal mm_interconnect_0_mm_reloj_0_avalon_slave_0_write                            : std_logic;                     -- mm_interconnect_0:mm_reloj_0_avalon_slave_0_write -> mm_reloj_0:write
	signal mm_interconnect_0_mm_reloj_0_avalon_slave_0_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:mm_reloj_0_avalon_slave_0_writedata -> mm_reloj_0:writedata
	signal mm_interconnect_0_new_sdram_controller_0_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	signal mm_interconnect_0_new_sdram_controller_0_s1_readdata                         : std_logic_vector(31 downto 0); -- new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	signal mm_interconnect_0_new_sdram_controller_0_s1_waitrequest                      : std_logic;                     -- new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	signal mm_interconnect_0_new_sdram_controller_0_s1_address                          : std_logic_vector(24 downto 0); -- mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	signal mm_interconnect_0_new_sdram_controller_0_s1_read                             : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_read -> mm_interconnect_0_new_sdram_controller_0_s1_read:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_byteenable                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> mm_interconnect_0_new_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid                    : std_logic;                     -- new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_0_new_sdram_controller_0_s1_write                            : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_write -> mm_interconnect_0_new_sdram_controller_0_s1_write:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	signal irq_mapper_receiver0_irq                                                     : std_logic;                     -- ps2_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                     : std_logic;                     -- mm_reloj_0:int_clk -> irq_mapper:receiver1_irq
	signal ensamblado_procesador_0_interrupt_receiver_irq                               : std_logic_vector(1 downto 0);  -- irq_mapper:sender_irq -> ensamblado_procesador_0:irq
	signal rst_controller_reset_out_reset                                               : std_logic;                     -- rst_controller:reset_out -> [ensamblado_procesador_0:reset, irq_mapper:reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:video_dma_controller_0_reset_reset_bridge_in_reset_reset, mm_reloj_0:Pcero, ps2_0:reset, sram_0:reset, video_dma_controller_0:reset, video_dual_clock_buffer_0:reset_stream_in, video_pll_0:ref_reset_reset]
	signal rst_controller_001_reset_out_reset                                           : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:new_sdram_controller_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal sys_sdram_pll_0_reset_source_reset                                           : std_logic;                     -- sys_sdram_pll_0:reset_source_reset -> rst_controller_001:reset_in0
	signal rst_controller_002_reset_out_reset                                           : std_logic;                     -- rst_controller_002:reset_out -> sys_sdram_pll_0:ref_reset_reset
	signal rst_controller_003_reset_out_reset                                           : std_logic;                     -- rst_controller_003:reset_out -> [video_dual_clock_buffer_0:reset_stream_out, video_vga_controller_0:reset]
	signal video_pll_0_reset_source_reset                                               : std_logic;                     -- video_pll_0:reset_source_reset -> rst_controller_003:reset_in0
	signal reset_reset_n_ports_inv                                                      : std_logic;                     -- reset_reset_n:inv -> [master_0:clk_reset_reset, rst_controller:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv                   : std_logic;                     -- mm_interconnect_0_new_sdram_controller_0_s1_read:inv -> new_sdram_controller_0:az_rd_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv             : std_logic_vector(3 downto 0);  -- mm_interconnect_0_new_sdram_controller_0_s1_byteenable:inv -> new_sdram_controller_0:az_be_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_new_sdram_controller_0_s1_write:inv -> new_sdram_controller_0:az_wr_n
	signal rst_controller_001_reset_out_reset_ports_inv                                 : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> new_sdram_controller_0:reset_n

begin

	ensamblado_procesador_0 : component ensamblado_procesador
		port map (
			reset         => rst_controller_reset_out_reset,                      --              reset.reset
			address       => ensamblado_procesador_0_avalon_master_address,       --      avalon_master.address
			writedata     => ensamblado_procesador_0_avalon_master_writedata,     --                   .writedata
			readdata      => ensamblado_procesador_0_avalon_master_readdata,      --                   .readdata
			read          => ensamblado_procesador_0_avalon_master_read,          --                   .read
			write         => ensamblado_procesador_0_avalon_master_write,         --                   .write
			byteenable    => ensamblado_procesador_0_avalon_master_byteenable,    --                   .byteenable
			waitrequest   => ensamblado_procesador_0_avalon_master_waitrequest,   --                   .waitrequest
			readdatavalid => ensamblado_procesador_0_avalon_master_readdatavalid, --                   .readdatavalid
			reloj         => sys_sdram_pll_0_sys_clk_clk,                         --         clock_sink.clk
			irq           => ensamblado_procesador_0_interrupt_receiver_irq,      -- interrupt_receiver.irq
			start         => start_bit                                            --        conduit_end.bit
		);

	master_0 : component disenyo_qsys_master_0
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => sys_sdram_pll_0_sys_clk_clk,   --          clk.clk
			clk_reset_reset      => reset_reset_n_ports_inv,       --    clk_reset.reset
			master_address       => master_0_master_address,       --       master.address
			master_readdata      => master_0_master_readdata,      --             .readdata
			master_read          => master_0_master_read,          --             .read
			master_write         => master_0_master_write,         --             .write
			master_writedata     => master_0_master_writedata,     --             .writedata
			master_waitrequest   => master_0_master_waitrequest,   --             .waitrequest
			master_readdatavalid => master_0_master_readdatavalid, --             .readdatavalid
			master_byteenable    => master_0_master_byteenable,    --             .byteenable
			master_reset_reset   => open                           -- master_reset.reset
		);

	mm_reloj_0 : component mm_reloj
		port map (
			read          => mm_interconnect_0_mm_reloj_0_avalon_slave_0_read,          --   avalon_slave_0.read
			write         => mm_interconnect_0_mm_reloj_0_avalon_slave_0_write,         --                 .write
			address       => mm_interconnect_0_mm_reloj_0_avalon_slave_0_address,       --                 .address
			writedata     => mm_interconnect_0_mm_reloj_0_avalon_slave_0_writedata,     --                 .writedata
			byteenable    => mm_interconnect_0_mm_reloj_0_avalon_slave_0_byteenable,    --                 .byteenable
			readdata      => mm_interconnect_0_mm_reloj_0_avalon_slave_0_readdata,      --                 .readdata
			waitrequest   => mm_interconnect_0_mm_reloj_0_avalon_slave_0_waitrequest,   --                 .waitrequest
			readdatavalid => mm_interconnect_0_mm_reloj_0_avalon_slave_0_readdatavalid, --                 .readdatavalid
			Pcero         => rst_controller_reset_out_reset,                            --       reset_sink.reset
			reloj         => sys_sdram_pll_0_sys_clk_clk,                               --       clock_sink.clk
			int_clk       => irq_mapper_receiver1_irq                                   -- interrupt_sender.irq
		);

	new_sdram_controller_0 : component disenyo_qsys_new_sdram_controller_0
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                      --   clk.clk
			reset_n        => rst_controller_001_reset_out_reset_ports_inv,                     -- reset.reset_n
			az_addr        => mm_interconnect_0_new_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_new_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_new_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_new_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_new_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                                  --  wire.export
			zs_ba          => sdram_wire_ba,                                                    --      .export
			zs_cas_n       => sdram_wire_cas_n,                                                 --      .export
			zs_cke         => sdram_wire_cke,                                                   --      .export
			zs_cs_n        => sdram_wire_cs_n,                                                  --      .export
			zs_dq          => sdram_wire_dq,                                                    --      .export
			zs_dqm         => sdram_wire_dqm,                                                   --      .export
			zs_ras_n       => sdram_wire_ras_n,                                                 --      .export
			zs_we_n        => sdram_wire_we_n                                                   --      .export
		);

	ps2_0 : component disenyo_qsys_ps2_0
		port map (
			clk         => sys_sdram_pll_0_sys_clk_clk,                          --                clk.clk
			reset       => rst_controller_reset_out_reset,                       --              reset.reset
			address     => mm_interconnect_0_ps2_0_avalon_ps2_slave_address(0),  --   avalon_ps2_slave.address
			chipselect  => mm_interconnect_0_ps2_0_avalon_ps2_slave_chipselect,  --                   .chipselect
			byteenable  => mm_interconnect_0_ps2_0_avalon_ps2_slave_byteenable,  --                   .byteenable
			read        => mm_interconnect_0_ps2_0_avalon_ps2_slave_read,        --                   .read
			write       => mm_interconnect_0_ps2_0_avalon_ps2_slave_write,       --                   .write
			writedata   => mm_interconnect_0_ps2_0_avalon_ps2_slave_writedata,   --                   .writedata
			readdata    => mm_interconnect_0_ps2_0_avalon_ps2_slave_readdata,    --                   .readdata
			waitrequest => mm_interconnect_0_ps2_0_avalon_ps2_slave_waitrequest, --                   .waitrequest
			irq         => irq_mapper_receiver0_irq,                             --          interrupt.irq
			PS2_CLK     => ps2_CLK,                                              -- external_interface.export
			PS2_DAT     => ps2_DAT                                               --                   .export
		);

	sram_0 : component disenyo_qsys_sram_0
		port map (
			clk           => sys_sdram_pll_0_sys_clk_clk,                              --                clk.clk
			reset         => rst_controller_reset_out_reset,                           --              reset.reset
			SRAM_DQ       => sram_DQ,                                                  -- external_interface.export
			SRAM_ADDR     => sram_ADDR,                                                --                   .export
			SRAM_LB_N     => sram_LB_N,                                                --                   .export
			SRAM_UB_N     => sram_UB_N,                                                --                   .export
			SRAM_CE_N     => sram_CE_N,                                                --                   .export
			SRAM_OE_N     => sram_OE_N,                                                --                   .export
			SRAM_WE_N     => sram_WE_N,                                                --                   .export
			address       => mm_interconnect_0_sram_0_avalon_sram_slave_address,       --  avalon_sram_slave.address
			byteenable    => mm_interconnect_0_sram_0_avalon_sram_slave_byteenable,    --                   .byteenable
			read          => mm_interconnect_0_sram_0_avalon_sram_slave_read,          --                   .read
			write         => mm_interconnect_0_sram_0_avalon_sram_slave_write,         --                   .write
			writedata     => mm_interconnect_0_sram_0_avalon_sram_slave_writedata,     --                   .writedata
			readdata      => mm_interconnect_0_sram_0_avalon_sram_slave_readdata,      --                   .readdata
			readdatavalid => mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid  --                   .readdatavalid
		);

	sys_sdram_pll_0 : component disenyo_qsys_sys_sdram_pll_0
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => rst_controller_002_reset_out_reset, --    ref_reset.reset
			sys_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                      --    sdram_clk.clk
			reset_source_reset => sys_sdram_pll_0_reset_source_reset  -- reset_source.reset
		);

	video_dma_controller_0 : component disenyo_qsys_video_dma_controller_0
		port map (
			clk                  => sys_sdram_pll_0_sys_clk_clk,                                                  --                      clk.clk
			reset                => rst_controller_reset_out_reset,                                               --                    reset.reset
			master_address       => video_dma_controller_0_avalon_dma_master_address,                             --        avalon_dma_master.address
			master_waitrequest   => video_dma_controller_0_avalon_dma_master_waitrequest,                         --                         .waitrequest
			master_arbiterlock   => video_dma_controller_0_avalon_dma_master_lock,                                --                         .lock
			master_read          => video_dma_controller_0_avalon_dma_master_read,                                --                         .read
			master_readdata      => video_dma_controller_0_avalon_dma_master_readdata,                            --                         .readdata
			master_readdatavalid => video_dma_controller_0_avalon_dma_master_readdatavalid,                       --                         .readdatavalid
			slave_address        => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_address,    -- avalon_dma_control_slave.address
			slave_byteenable     => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_byteenable, --                         .byteenable
			slave_read           => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_read,       --                         .read
			slave_write          => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_write,      --                         .write
			slave_writedata      => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_writedata,  --                         .writedata
			slave_readdata       => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_readdata,   --                         .readdata
			stream_ready         => video_dma_controller_0_avalon_pixel_source_ready,                             --      avalon_pixel_source.ready
			stream_data          => video_dma_controller_0_avalon_pixel_source_data,                              --                         .data
			stream_startofpacket => video_dma_controller_0_avalon_pixel_source_startofpacket,                     --                         .startofpacket
			stream_endofpacket   => video_dma_controller_0_avalon_pixel_source_endofpacket,                       --                         .endofpacket
			stream_valid         => video_dma_controller_0_avalon_pixel_source_valid                              --                         .valid
		);

	video_dual_clock_buffer_0 : component disenyo_qsys_video_dual_clock_buffer_0
		port map (
			clk_stream_in            => sys_sdram_pll_0_sys_clk_clk,                                     --         clock_stream_in.clk
			reset_stream_in          => rst_controller_reset_out_reset,                                  --         reset_stream_in.reset
			clk_stream_out           => video_pll_0_vga_clk_clk,                                         --        clock_stream_out.clk
			reset_stream_out         => rst_controller_003_reset_out_reset,                              --        reset_stream_out.reset
			stream_in_ready          => video_dma_controller_0_avalon_pixel_source_ready,                --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => video_dma_controller_0_avalon_pixel_source_startofpacket,        --                        .startofpacket
			stream_in_endofpacket    => video_dma_controller_0_avalon_pixel_source_endofpacket,          --                        .endofpacket
			stream_in_valid          => video_dma_controller_0_avalon_pixel_source_valid,                --                        .valid
			stream_in_data           => video_dma_controller_0_avalon_pixel_source_data,                 --                        .data
			stream_out_ready         => video_dual_clock_buffer_0_avalon_dc_buffer_source_ready,         -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket, --                        .startofpacket
			stream_out_endofpacket   => video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket,   --                        .endofpacket
			stream_out_valid         => video_dual_clock_buffer_0_avalon_dc_buffer_source_valid,         --                        .valid
			stream_out_data          => video_dual_clock_buffer_0_avalon_dc_buffer_source_data           --                        .data
		);

	video_pll_0 : component disenyo_qsys_video_pll_0
		port map (
			ref_clk_clk        => sys_sdram_pll_0_sys_clk_clk,    --      ref_clk.clk
			ref_reset_reset    => rst_controller_reset_out_reset, --    ref_reset.reset
			vga_clk_clk        => video_pll_0_vga_clk_clk,        --      vga_clk.clk
			reset_source_reset => video_pll_0_reset_source_reset  -- reset_source.reset
		);

	video_vga_controller_0 : component disenyo_qsys_video_vga_controller_0
		port map (
			clk           => video_pll_0_vga_clk_clk,                                         --                clk.clk
			reset         => rst_controller_003_reset_out_reset,                              --              reset.reset
			data          => video_dual_clock_buffer_0_avalon_dc_buffer_source_data,          --    avalon_vga_sink.data
			startofpacket => video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket, --                   .startofpacket
			endofpacket   => video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket,   --                   .endofpacket
			valid         => video_dual_clock_buffer_0_avalon_dc_buffer_source_valid,         --                   .valid
			ready         => video_dual_clock_buffer_0_avalon_dc_buffer_source_ready,         --                   .ready
			VGA_CLK       => vga_CLK,                                                         -- external_interface.export
			VGA_HS        => vga_HS,                                                          --                   .export
			VGA_VS        => vga_VS,                                                          --                   .export
			VGA_BLANK     => vga_BLANK,                                                       --                   .export
			VGA_SYNC      => vga_SYNC,                                                        --                   .export
			VGA_R         => vga_R,                                                           --                   .export
			VGA_G         => vga_G,                                                           --                   .export
			VGA_B         => vga_B                                                            --                   .export
		);

	mm_interconnect_0 : component disenyo_qsys_mm_interconnect_0
		port map (
			sys_sdram_pll_0_sys_clk_clk                                => sys_sdram_pll_0_sys_clk_clk,                                                  --                            sys_sdram_pll_0_sys_clk.clk
			master_0_clk_reset_reset_bridge_in_reset_reset             => rst_controller_reset_out_reset,                                               --           master_0_clk_reset_reset_bridge_in_reset.reset
			new_sdram_controller_0_reset_reset_bridge_in_reset_reset   => rst_controller_001_reset_out_reset,                                           -- new_sdram_controller_0_reset_reset_bridge_in_reset.reset
			video_dma_controller_0_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                                               -- video_dma_controller_0_reset_reset_bridge_in_reset.reset
			ensamblado_procesador_0_avalon_master_address              => ensamblado_procesador_0_avalon_master_address,                                --              ensamblado_procesador_0_avalon_master.address
			ensamblado_procesador_0_avalon_master_waitrequest          => ensamblado_procesador_0_avalon_master_waitrequest,                            --                                                   .waitrequest
			ensamblado_procesador_0_avalon_master_byteenable           => ensamblado_procesador_0_avalon_master_byteenable,                             --                                                   .byteenable
			ensamblado_procesador_0_avalon_master_read                 => ensamblado_procesador_0_avalon_master_read,                                   --                                                   .read
			ensamblado_procesador_0_avalon_master_readdata             => ensamblado_procesador_0_avalon_master_readdata,                               --                                                   .readdata
			ensamblado_procesador_0_avalon_master_readdatavalid        => ensamblado_procesador_0_avalon_master_readdatavalid,                          --                                                   .readdatavalid
			ensamblado_procesador_0_avalon_master_write                => ensamblado_procesador_0_avalon_master_write,                                  --                                                   .write
			ensamblado_procesador_0_avalon_master_writedata            => ensamblado_procesador_0_avalon_master_writedata,                              --                                                   .writedata
			master_0_master_address                                    => master_0_master_address,                                                      --                                    master_0_master.address
			master_0_master_waitrequest                                => master_0_master_waitrequest,                                                  --                                                   .waitrequest
			master_0_master_byteenable                                 => master_0_master_byteenable,                                                   --                                                   .byteenable
			master_0_master_read                                       => master_0_master_read,                                                         --                                                   .read
			master_0_master_readdata                                   => master_0_master_readdata,                                                     --                                                   .readdata
			master_0_master_readdatavalid                              => master_0_master_readdatavalid,                                                --                                                   .readdatavalid
			master_0_master_write                                      => master_0_master_write,                                                        --                                                   .write
			master_0_master_writedata                                  => master_0_master_writedata,                                                    --                                                   .writedata
			video_dma_controller_0_avalon_dma_master_address           => video_dma_controller_0_avalon_dma_master_address,                             --           video_dma_controller_0_avalon_dma_master.address
			video_dma_controller_0_avalon_dma_master_waitrequest       => video_dma_controller_0_avalon_dma_master_waitrequest,                         --                                                   .waitrequest
			video_dma_controller_0_avalon_dma_master_read              => video_dma_controller_0_avalon_dma_master_read,                                --                                                   .read
			video_dma_controller_0_avalon_dma_master_readdata          => video_dma_controller_0_avalon_dma_master_readdata,                            --                                                   .readdata
			video_dma_controller_0_avalon_dma_master_readdatavalid     => video_dma_controller_0_avalon_dma_master_readdatavalid,                       --                                                   .readdatavalid
			video_dma_controller_0_avalon_dma_master_lock              => video_dma_controller_0_avalon_dma_master_lock,                                --                                                   .lock
			mm_reloj_0_avalon_slave_0_address                          => mm_interconnect_0_mm_reloj_0_avalon_slave_0_address,                          --                          mm_reloj_0_avalon_slave_0.address
			mm_reloj_0_avalon_slave_0_write                            => mm_interconnect_0_mm_reloj_0_avalon_slave_0_write,                            --                                                   .write
			mm_reloj_0_avalon_slave_0_read                             => mm_interconnect_0_mm_reloj_0_avalon_slave_0_read,                             --                                                   .read
			mm_reloj_0_avalon_slave_0_readdata                         => mm_interconnect_0_mm_reloj_0_avalon_slave_0_readdata,                         --                                                   .readdata
			mm_reloj_0_avalon_slave_0_writedata                        => mm_interconnect_0_mm_reloj_0_avalon_slave_0_writedata,                        --                                                   .writedata
			mm_reloj_0_avalon_slave_0_byteenable                       => mm_interconnect_0_mm_reloj_0_avalon_slave_0_byteenable,                       --                                                   .byteenable
			mm_reloj_0_avalon_slave_0_readdatavalid                    => mm_interconnect_0_mm_reloj_0_avalon_slave_0_readdatavalid,                    --                                                   .readdatavalid
			mm_reloj_0_avalon_slave_0_waitrequest                      => mm_interconnect_0_mm_reloj_0_avalon_slave_0_waitrequest,                      --                                                   .waitrequest
			new_sdram_controller_0_s1_address                          => mm_interconnect_0_new_sdram_controller_0_s1_address,                          --                          new_sdram_controller_0_s1.address
			new_sdram_controller_0_s1_write                            => mm_interconnect_0_new_sdram_controller_0_s1_write,                            --                                                   .write
			new_sdram_controller_0_s1_read                             => mm_interconnect_0_new_sdram_controller_0_s1_read,                             --                                                   .read
			new_sdram_controller_0_s1_readdata                         => mm_interconnect_0_new_sdram_controller_0_s1_readdata,                         --                                                   .readdata
			new_sdram_controller_0_s1_writedata                        => mm_interconnect_0_new_sdram_controller_0_s1_writedata,                        --                                                   .writedata
			new_sdram_controller_0_s1_byteenable                       => mm_interconnect_0_new_sdram_controller_0_s1_byteenable,                       --                                                   .byteenable
			new_sdram_controller_0_s1_readdatavalid                    => mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid,                    --                                                   .readdatavalid
			new_sdram_controller_0_s1_waitrequest                      => mm_interconnect_0_new_sdram_controller_0_s1_waitrequest,                      --                                                   .waitrequest
			new_sdram_controller_0_s1_chipselect                       => mm_interconnect_0_new_sdram_controller_0_s1_chipselect,                       --                                                   .chipselect
			ps2_0_avalon_ps2_slave_address                             => mm_interconnect_0_ps2_0_avalon_ps2_slave_address,                             --                             ps2_0_avalon_ps2_slave.address
			ps2_0_avalon_ps2_slave_write                               => mm_interconnect_0_ps2_0_avalon_ps2_slave_write,                               --                                                   .write
			ps2_0_avalon_ps2_slave_read                                => mm_interconnect_0_ps2_0_avalon_ps2_slave_read,                                --                                                   .read
			ps2_0_avalon_ps2_slave_readdata                            => mm_interconnect_0_ps2_0_avalon_ps2_slave_readdata,                            --                                                   .readdata
			ps2_0_avalon_ps2_slave_writedata                           => mm_interconnect_0_ps2_0_avalon_ps2_slave_writedata,                           --                                                   .writedata
			ps2_0_avalon_ps2_slave_byteenable                          => mm_interconnect_0_ps2_0_avalon_ps2_slave_byteenable,                          --                                                   .byteenable
			ps2_0_avalon_ps2_slave_waitrequest                         => mm_interconnect_0_ps2_0_avalon_ps2_slave_waitrequest,                         --                                                   .waitrequest
			ps2_0_avalon_ps2_slave_chipselect                          => mm_interconnect_0_ps2_0_avalon_ps2_slave_chipselect,                          --                                                   .chipselect
			sram_0_avalon_sram_slave_address                           => mm_interconnect_0_sram_0_avalon_sram_slave_address,                           --                           sram_0_avalon_sram_slave.address
			sram_0_avalon_sram_slave_write                             => mm_interconnect_0_sram_0_avalon_sram_slave_write,                             --                                                   .write
			sram_0_avalon_sram_slave_read                              => mm_interconnect_0_sram_0_avalon_sram_slave_read,                              --                                                   .read
			sram_0_avalon_sram_slave_readdata                          => mm_interconnect_0_sram_0_avalon_sram_slave_readdata,                          --                                                   .readdata
			sram_0_avalon_sram_slave_writedata                         => mm_interconnect_0_sram_0_avalon_sram_slave_writedata,                         --                                                   .writedata
			sram_0_avalon_sram_slave_byteenable                        => mm_interconnect_0_sram_0_avalon_sram_slave_byteenable,                        --                                                   .byteenable
			sram_0_avalon_sram_slave_readdatavalid                     => mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid,                     --                                                   .readdatavalid
			video_dma_controller_0_avalon_dma_control_slave_address    => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_address,    --    video_dma_controller_0_avalon_dma_control_slave.address
			video_dma_controller_0_avalon_dma_control_slave_write      => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_write,      --                                                   .write
			video_dma_controller_0_avalon_dma_control_slave_read       => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_read,       --                                                   .read
			video_dma_controller_0_avalon_dma_control_slave_readdata   => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_readdata,   --                                                   .readdata
			video_dma_controller_0_avalon_dma_control_slave_writedata  => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_writedata,  --                                                   .writedata
			video_dma_controller_0_avalon_dma_control_slave_byteenable => mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_byteenable  --                                                   .byteenable
		);

	irq_mapper : component disenyo_qsys_irq_mapper
		port map (
			clk           => sys_sdram_pll_0_sys_clk_clk,                    --       clk.clk
			reset         => rst_controller_reset_out_reset,                 -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,                       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,                       -- receiver1.irq
			sender_irq    => ensamblado_procesador_0_interrupt_receiver_irq  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,    --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_sdram_pll_0_reset_source_reset, -- reset_in0.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => video_pll_0_reset_source_reset,     -- reset_in0.reset
			clk            => video_pll_0_vga_clk_clk,            --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_read;

	mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_byteenable;

	mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of disenyo_qsys
