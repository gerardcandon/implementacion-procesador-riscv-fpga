-- disenyo_qsys.vhd

-- Generated using ACDS version 19.1 670

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity disenyo_qsys is
	port (
		clk_clk          : in    std_logic                     := '0';             --        clk.clk
		reset_reset_n    : in    std_logic                     := '0';             --      reset.reset_n
		sdram_clk_clk    : out   std_logic;                                        --  sdram_clk.clk
		sdram_wire_addr  : out   std_logic_vector(12 downto 0);                    -- sdram_wire.addr
		sdram_wire_ba    : out   std_logic_vector(1 downto 0);                     --           .ba
		sdram_wire_cas_n : out   std_logic;                                        --           .cas_n
		sdram_wire_cke   : out   std_logic;                                        --           .cke
		sdram_wire_cs_n  : out   std_logic;                                        --           .cs_n
		sdram_wire_dq    : inout std_logic_vector(31 downto 0) := (others => '0'); --           .dq
		sdram_wire_dqm   : out   std_logic_vector(3 downto 0);                     --           .dqm
		sdram_wire_ras_n : out   std_logic;                                        --           .ras_n
		sdram_wire_we_n  : out   std_logic                                         --           .we_n
	);
end entity disenyo_qsys;

architecture rtl of disenyo_qsys is
	component ensamblado_procesador is
		port (
			reloj           : in  std_logic                     := 'X';             -- clk
			Pcero           : in  std_logic                     := 'X';             -- reset
			address_M       : out std_logic_vector(31 downto 0);                    -- address
			byteenable_M    : out std_logic_vector(3 downto 0);                     -- byteenable
			read_M          : out std_logic;                                        -- read
			readdata_M      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			readdatavalid_M : in  std_logic                     := 'X';             -- readdatavalid
			waitrequest_M   : in  std_logic                     := 'X';             -- waitrequest
			write_M         : out std_logic;                                        -- write
			writedata_M     : out std_logic_vector(31 downto 0);                    -- writedata
			address_B       : out std_logic_vector(31 downto 0);                    -- address
			readdata_B      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			read_B          : out std_logic;                                        -- read
			byteenable_B    : out std_logic_vector(3 downto 0);                     -- byteenable
			waitrequest_B   : in  std_logic                     := 'X';             -- waitrequest
			readdatavalid_B : in  std_logic                     := 'X'              -- readdatavalid
		);
	end component ensamblado_procesador;

	component disenyo_qsys_master_0 is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component disenyo_qsys_master_0;

	component disenyo_qsys_new_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component disenyo_qsys_new_sdram_controller_0;

	component disenyo_qsys_sys_sdram_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component disenyo_qsys_sys_sdram_pll_0;

	component disenyo_qsys_mm_interconnect_0 is
		port (
			sys_sdram_pll_0_sys_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			ensamblado_procesador_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			master_0_clk_reset_reset_bridge_in_reset_reset                 : in  std_logic                     := 'X';             -- reset
			ensamblado_procesador_0_avalon_master_B_address                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			ensamblado_procesador_0_avalon_master_B_waitrequest            : out std_logic;                                        -- waitrequest
			ensamblado_procesador_0_avalon_master_B_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ensamblado_procesador_0_avalon_master_B_read                   : in  std_logic                     := 'X';             -- read
			ensamblado_procesador_0_avalon_master_B_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			ensamblado_procesador_0_avalon_master_B_readdatavalid          : out std_logic;                                        -- readdatavalid
			ensamblado_procesador_0_avalon_master_M_address                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			ensamblado_procesador_0_avalon_master_M_waitrequest            : out std_logic;                                        -- waitrequest
			ensamblado_procesador_0_avalon_master_M_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ensamblado_procesador_0_avalon_master_M_read                   : in  std_logic                     := 'X';             -- read
			ensamblado_procesador_0_avalon_master_M_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			ensamblado_procesador_0_avalon_master_M_readdatavalid          : out std_logic;                                        -- readdatavalid
			ensamblado_procesador_0_avalon_master_M_write                  : in  std_logic                     := 'X';             -- write
			ensamblado_procesador_0_avalon_master_M_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			master_0_master_address                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			master_0_master_waitrequest                                    : out std_logic;                                        -- waitrequest
			master_0_master_byteenable                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			master_0_master_read                                           : in  std_logic                     := 'X';             -- read
			master_0_master_readdata                                       : out std_logic_vector(31 downto 0);                    -- readdata
			master_0_master_readdatavalid                                  : out std_logic;                                        -- readdatavalid
			master_0_master_write                                          : in  std_logic                     := 'X';             -- write
			master_0_master_writedata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			new_sdram_controller_0_s1_address                              : out std_logic_vector(24 downto 0);                    -- address
			new_sdram_controller_0_s1_write                                : out std_logic;                                        -- write
			new_sdram_controller_0_s1_read                                 : out std_logic;                                        -- read
			new_sdram_controller_0_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			new_sdram_controller_0_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			new_sdram_controller_0_s1_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			new_sdram_controller_0_s1_readdatavalid                        : in  std_logic                     := 'X';             -- readdatavalid
			new_sdram_controller_0_s1_waitrequest                          : in  std_logic                     := 'X';             -- waitrequest
			new_sdram_controller_0_s1_chipselect                           : out std_logic                                         -- chipselect
		);
	end component disenyo_qsys_mm_interconnect_0;

	component disenyo_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			reset_in2      : in  std_logic := 'X'; -- reset_in2.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component disenyo_qsys_rst_controller;

	component disenyo_qsys_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component disenyo_qsys_rst_controller_002;

	signal sys_sdram_pll_0_sys_clk_clk                                      : std_logic;                     -- sys_sdram_pll_0:sys_clk_clk -> [ensamblado_procesador_0:reloj, master_0:clk_clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, new_sdram_controller_0:clk, rst_controller:clk]
	signal ensamblado_procesador_0_avalon_master_b_readdata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:ensamblado_procesador_0_avalon_master_B_readdata -> ensamblado_procesador_0:readdata_B
	signal ensamblado_procesador_0_avalon_master_b_waitrequest              : std_logic;                     -- mm_interconnect_0:ensamblado_procesador_0_avalon_master_B_waitrequest -> ensamblado_procesador_0:waitrequest_B
	signal ensamblado_procesador_0_avalon_master_b_address                  : std_logic_vector(31 downto 0); -- ensamblado_procesador_0:address_B -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_B_address
	signal ensamblado_procesador_0_avalon_master_b_read                     : std_logic;                     -- ensamblado_procesador_0:read_B -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_B_read
	signal ensamblado_procesador_0_avalon_master_b_byteenable               : std_logic_vector(3 downto 0);  -- ensamblado_procesador_0:byteenable_B -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_B_byteenable
	signal ensamblado_procesador_0_avalon_master_b_readdatavalid            : std_logic;                     -- mm_interconnect_0:ensamblado_procesador_0_avalon_master_B_readdatavalid -> ensamblado_procesador_0:readdatavalid_B
	signal ensamblado_procesador_0_avalon_master_m_readdata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:ensamblado_procesador_0_avalon_master_M_readdata -> ensamblado_procesador_0:readdata_M
	signal ensamblado_procesador_0_avalon_master_m_waitrequest              : std_logic;                     -- mm_interconnect_0:ensamblado_procesador_0_avalon_master_M_waitrequest -> ensamblado_procesador_0:waitrequest_M
	signal ensamblado_procesador_0_avalon_master_m_address                  : std_logic_vector(31 downto 0); -- ensamblado_procesador_0:address_M -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_M_address
	signal ensamblado_procesador_0_avalon_master_m_byteenable               : std_logic_vector(3 downto 0);  -- ensamblado_procesador_0:byteenable_M -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_M_byteenable
	signal ensamblado_procesador_0_avalon_master_m_read                     : std_logic;                     -- ensamblado_procesador_0:read_M -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_M_read
	signal ensamblado_procesador_0_avalon_master_m_readdatavalid            : std_logic;                     -- mm_interconnect_0:ensamblado_procesador_0_avalon_master_M_readdatavalid -> ensamblado_procesador_0:readdatavalid_M
	signal ensamblado_procesador_0_avalon_master_m_write                    : std_logic;                     -- ensamblado_procesador_0:write_M -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_M_write
	signal ensamblado_procesador_0_avalon_master_m_writedata                : std_logic_vector(31 downto 0); -- ensamblado_procesador_0:writedata_M -> mm_interconnect_0:ensamblado_procesador_0_avalon_master_M_writedata
	signal master_0_master_readdata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	signal master_0_master_waitrequest                                      : std_logic;                     -- mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	signal master_0_master_address                                          : std_logic_vector(31 downto 0); -- master_0:master_address -> mm_interconnect_0:master_0_master_address
	signal master_0_master_read                                             : std_logic;                     -- master_0:master_read -> mm_interconnect_0:master_0_master_read
	signal master_0_master_byteenable                                       : std_logic_vector(3 downto 0);  -- master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	signal master_0_master_readdatavalid                                    : std_logic;                     -- mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	signal master_0_master_write                                            : std_logic;                     -- master_0:master_write -> mm_interconnect_0:master_0_master_write
	signal master_0_master_writedata                                        : std_logic_vector(31 downto 0); -- master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	signal mm_interconnect_0_new_sdram_controller_0_s1_chipselect           : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	signal mm_interconnect_0_new_sdram_controller_0_s1_readdata             : std_logic_vector(31 downto 0); -- new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	signal mm_interconnect_0_new_sdram_controller_0_s1_waitrequest          : std_logic;                     -- new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	signal mm_interconnect_0_new_sdram_controller_0_s1_address              : std_logic_vector(24 downto 0); -- mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	signal mm_interconnect_0_new_sdram_controller_0_s1_read                 : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_read -> mm_interconnect_0_new_sdram_controller_0_s1_read:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> mm_interconnect_0_new_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid        : std_logic;                     -- new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_0_new_sdram_controller_0_s1_write                : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_write -> mm_interconnect_0_new_sdram_controller_0_s1_write:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	signal rst_controller_reset_out_reset                                   : std_logic;                     -- rst_controller:reset_out -> [ensamblado_procesador_0:Pcero, mm_interconnect_0:ensamblado_procesador_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal master_0_master_reset_reset                                      : std_logic;                     -- master_0:master_reset_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal sys_sdram_pll_0_reset_source_reset                               : std_logic;                     -- sys_sdram_pll_0:reset_source_reset -> [rst_controller:reset_in2, rst_controller_001:reset_in2]
	signal rst_controller_001_reset_out_reset                               : std_logic;                     -- rst_controller_001:reset_out -> master_0:clk_reset_reset
	signal rst_controller_002_reset_out_reset                               : std_logic;                     -- rst_controller_002:reset_out -> sys_sdram_pll_0:ref_reset_reset
	signal reset_reset_n_ports_inv                                          : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv       : std_logic;                     -- mm_interconnect_0_new_sdram_controller_0_s1_read:inv -> new_sdram_controller_0:az_rd_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv : std_logic_vector(3 downto 0);  -- mm_interconnect_0_new_sdram_controller_0_s1_byteenable:inv -> new_sdram_controller_0:az_be_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv      : std_logic;                     -- mm_interconnect_0_new_sdram_controller_0_s1_write:inv -> new_sdram_controller_0:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                         : std_logic;                     -- rst_controller_reset_out_reset:inv -> new_sdram_controller_0:reset_n

begin

	ensamblado_procesador_0 : component ensamblado_procesador
		port map (
			reloj           => sys_sdram_pll_0_sys_clk_clk,                           --      clock_sink.clk
			Pcero           => rst_controller_reset_out_reset,                        --      reset_sink.reset
			address_M       => ensamblado_procesador_0_avalon_master_m_address,       -- avalon_master_M.address
			byteenable_M    => ensamblado_procesador_0_avalon_master_m_byteenable,    --                .byteenable
			read_M          => ensamblado_procesador_0_avalon_master_m_read,          --                .read
			readdata_M      => ensamblado_procesador_0_avalon_master_m_readdata,      --                .readdata
			readdatavalid_M => ensamblado_procesador_0_avalon_master_m_readdatavalid, --                .readdatavalid
			waitrequest_M   => ensamblado_procesador_0_avalon_master_m_waitrequest,   --                .waitrequest
			write_M         => ensamblado_procesador_0_avalon_master_m_write,         --                .write
			writedata_M     => ensamblado_procesador_0_avalon_master_m_writedata,     --                .writedata
			address_B       => ensamblado_procesador_0_avalon_master_b_address,       -- avalon_master_B.address
			readdata_B      => ensamblado_procesador_0_avalon_master_b_readdata,      --                .readdata
			read_B          => ensamblado_procesador_0_avalon_master_b_read,          --                .read
			byteenable_B    => ensamblado_procesador_0_avalon_master_b_byteenable,    --                .byteenable
			waitrequest_B   => ensamblado_procesador_0_avalon_master_b_waitrequest,   --                .waitrequest
			readdatavalid_B => ensamblado_procesador_0_avalon_master_b_readdatavalid  --                .readdatavalid
		);

	master_0 : component disenyo_qsys_master_0
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => sys_sdram_pll_0_sys_clk_clk,        --          clk.clk
			clk_reset_reset      => rst_controller_001_reset_out_reset, --    clk_reset.reset
			master_address       => master_0_master_address,            --       master.address
			master_readdata      => master_0_master_readdata,           --             .readdata
			master_read          => master_0_master_read,               --             .read
			master_write         => master_0_master_write,              --             .write
			master_writedata     => master_0_master_writedata,          --             .writedata
			master_waitrequest   => master_0_master_waitrequest,        --             .waitrequest
			master_readdatavalid => master_0_master_readdatavalid,      --             .readdatavalid
			master_byteenable    => master_0_master_byteenable,         --             .byteenable
			master_reset_reset   => master_0_master_reset_reset         -- master_reset.reset
		);

	new_sdram_controller_0 : component disenyo_qsys_new_sdram_controller_0
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                      --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                         -- reset.reset_n
			az_addr        => mm_interconnect_0_new_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_new_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_new_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_new_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_new_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                                  --  wire.export
			zs_ba          => sdram_wire_ba,                                                    --      .export
			zs_cas_n       => sdram_wire_cas_n,                                                 --      .export
			zs_cke         => sdram_wire_cke,                                                   --      .export
			zs_cs_n        => sdram_wire_cs_n,                                                  --      .export
			zs_dq          => sdram_wire_dq,                                                    --      .export
			zs_dqm         => sdram_wire_dqm,                                                   --      .export
			zs_ras_n       => sdram_wire_ras_n,                                                 --      .export
			zs_we_n        => sdram_wire_we_n                                                   --      .export
		);

	sys_sdram_pll_0 : component disenyo_qsys_sys_sdram_pll_0
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => rst_controller_002_reset_out_reset, --    ref_reset.reset
			sys_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                      --    sdram_clk.clk
			reset_source_reset => sys_sdram_pll_0_reset_source_reset  -- reset_source.reset
		);

	mm_interconnect_0 : component disenyo_qsys_mm_interconnect_0
		port map (
			sys_sdram_pll_0_sys_clk_clk                                    => sys_sdram_pll_0_sys_clk_clk,                               --                                  sys_sdram_pll_0_sys_clk.clk
			ensamblado_procesador_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- ensamblado_procesador_0_reset_sink_reset_bridge_in_reset.reset
			master_0_clk_reset_reset_bridge_in_reset_reset                 => rst_controller_reset_out_reset,                            --                 master_0_clk_reset_reset_bridge_in_reset.reset
			ensamblado_procesador_0_avalon_master_B_address                => ensamblado_procesador_0_avalon_master_b_address,           --                  ensamblado_procesador_0_avalon_master_B.address
			ensamblado_procesador_0_avalon_master_B_waitrequest            => ensamblado_procesador_0_avalon_master_b_waitrequest,       --                                                         .waitrequest
			ensamblado_procesador_0_avalon_master_B_byteenable             => ensamblado_procesador_0_avalon_master_b_byteenable,        --                                                         .byteenable
			ensamblado_procesador_0_avalon_master_B_read                   => ensamblado_procesador_0_avalon_master_b_read,              --                                                         .read
			ensamblado_procesador_0_avalon_master_B_readdata               => ensamblado_procesador_0_avalon_master_b_readdata,          --                                                         .readdata
			ensamblado_procesador_0_avalon_master_B_readdatavalid          => ensamblado_procesador_0_avalon_master_b_readdatavalid,     --                                                         .readdatavalid
			ensamblado_procesador_0_avalon_master_M_address                => ensamblado_procesador_0_avalon_master_m_address,           --                  ensamblado_procesador_0_avalon_master_M.address
			ensamblado_procesador_0_avalon_master_M_waitrequest            => ensamblado_procesador_0_avalon_master_m_waitrequest,       --                                                         .waitrequest
			ensamblado_procesador_0_avalon_master_M_byteenable             => ensamblado_procesador_0_avalon_master_m_byteenable,        --                                                         .byteenable
			ensamblado_procesador_0_avalon_master_M_read                   => ensamblado_procesador_0_avalon_master_m_read,              --                                                         .read
			ensamblado_procesador_0_avalon_master_M_readdata               => ensamblado_procesador_0_avalon_master_m_readdata,          --                                                         .readdata
			ensamblado_procesador_0_avalon_master_M_readdatavalid          => ensamblado_procesador_0_avalon_master_m_readdatavalid,     --                                                         .readdatavalid
			ensamblado_procesador_0_avalon_master_M_write                  => ensamblado_procesador_0_avalon_master_m_write,             --                                                         .write
			ensamblado_procesador_0_avalon_master_M_writedata              => ensamblado_procesador_0_avalon_master_m_writedata,         --                                                         .writedata
			master_0_master_address                                        => master_0_master_address,                                   --                                          master_0_master.address
			master_0_master_waitrequest                                    => master_0_master_waitrequest,                               --                                                         .waitrequest
			master_0_master_byteenable                                     => master_0_master_byteenable,                                --                                                         .byteenable
			master_0_master_read                                           => master_0_master_read,                                      --                                                         .read
			master_0_master_readdata                                       => master_0_master_readdata,                                  --                                                         .readdata
			master_0_master_readdatavalid                                  => master_0_master_readdatavalid,                             --                                                         .readdatavalid
			master_0_master_write                                          => master_0_master_write,                                     --                                                         .write
			master_0_master_writedata                                      => master_0_master_writedata,                                 --                                                         .writedata
			new_sdram_controller_0_s1_address                              => mm_interconnect_0_new_sdram_controller_0_s1_address,       --                                new_sdram_controller_0_s1.address
			new_sdram_controller_0_s1_write                                => mm_interconnect_0_new_sdram_controller_0_s1_write,         --                                                         .write
			new_sdram_controller_0_s1_read                                 => mm_interconnect_0_new_sdram_controller_0_s1_read,          --                                                         .read
			new_sdram_controller_0_s1_readdata                             => mm_interconnect_0_new_sdram_controller_0_s1_readdata,      --                                                         .readdata
			new_sdram_controller_0_s1_writedata                            => mm_interconnect_0_new_sdram_controller_0_s1_writedata,     --                                                         .writedata
			new_sdram_controller_0_s1_byteenable                           => mm_interconnect_0_new_sdram_controller_0_s1_byteenable,    --                                                         .byteenable
			new_sdram_controller_0_s1_readdatavalid                        => mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid, --                                                         .readdatavalid
			new_sdram_controller_0_s1_waitrequest                          => mm_interconnect_0_new_sdram_controller_0_s1_waitrequest,   --                                                         .waitrequest
			new_sdram_controller_0_s1_chipselect                           => mm_interconnect_0_new_sdram_controller_0_s1_chipselect     --                                                         .chipselect
		);

	rst_controller : component disenyo_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => master_0_master_reset_reset,        -- reset_in1.reset
			reset_in2      => sys_sdram_pll_0_reset_source_reset, -- reset_in2.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component disenyo_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => master_0_master_reset_reset,        -- reset_in1.reset
			reset_in2      => sys_sdram_pll_0_reset_source_reset, -- reset_in2.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component disenyo_qsys_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_read;

	mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_byteenable;

	mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of disenyo_qsys
