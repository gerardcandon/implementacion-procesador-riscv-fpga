-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions and other 
-- software and tools, and its AMPP partner logic functions, and any output 
-- files from any of the foregoing (including device programming or simulation 
-- files), and any associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License Subscription 
-- Agreement, Intel FPGA IP License Agreement, or other applicable 
-- license agreement, including, without limitation, that your use is for the 
-- sole purpose of programming logic devices manufactured by Intel and sold by 
-- Intel or its authorized distributors.  Please refer to the applicable 
-- agreement for further details.


-- $Id: //acds/main/ip/sopc/components/verification/altera_tristate_conduit_bfm/altera_tristate_conduit_bfm.sv.terp#7 $
-- $Revision: #7 $
-- $Date: 2010/08/05 $
-- $Author: klong $
-------------------------------------------------------------------------------
-- =head1 NAME
-- altera_conduit_bfm
-- =head1 SYNOPSIS
-- Bus Functional Model (BFM) for a Standard Conduit BFM
-------------------------------------------------------------------------------
-- =head1 DESCRIPTION
-- This is a Bus Functional Model (BFM) VHDL package for a Standard Conduit Master.
-- This package provides the API that will be used to get the value of the sampled
-- input/bidirection port or set the value to be driven to the output ports.
-- This BFM's HDL is been generated through terp file in Qsys/SOPC Builder.
-- Generation parameters:
-- output_name:                  altera_conduit_bfm
-- role:width:direction:         CLK:1:bidir,DAT:1:bidir
-- clocked                       0
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.all;



package altera_conduit_bfm_vhdl_pkg is

   -- output signal register
   type altera_conduit_bfm_out_trans_t is record
      sig_CLK_out     : std_logic_vector(0 downto 0);
      sig_CLK_oe      : std_logic;
      sig_DAT_out     : std_logic_vector(0 downto 0);
      sig_DAT_oe      : std_logic;
   end record;
   
   shared variable out_trans        : altera_conduit_bfm_out_trans_t;

   -- input signal register
   signal sig_CLK_in      : std_logic_vector(0 downto 0);
   signal sig_DAT_in      : std_logic_vector(0 downto 0);

   -- VHDL Procedure API
   
   -- get CLK value
   procedure get_CLK             (signal_value : out std_logic_vector(0 downto 0));
   
   -- set CLK value
   procedure set_CLK             (signal_value : in std_logic_vector(0 downto 0));
   
   -- set CLK input / output direction
   procedure set_CLK_oe          (signal_value : in std_logic);
   
   -- get DAT value
   procedure get_DAT             (signal_value : out std_logic_vector(0 downto 0));
   
   -- set DAT value
   procedure set_DAT             (signal_value : in std_logic_vector(0 downto 0));
   
   -- set DAT input / output direction
   procedure set_DAT_oe          (signal_value : in std_logic);
   
   -- VHDL Event API

   procedure event_CLK_change;   

   procedure event_DAT_change;   

end altera_conduit_bfm_vhdl_pkg;

package body altera_conduit_bfm_vhdl_pkg is
   
   procedure get_CLK             (signal_value : out std_logic_vector(0 downto 0)) is
   begin

      signal_value := sig_CLK_in;
   
   end procedure get_CLK;
   
   procedure set_CLK             (signal_value : in std_logic_vector(0 downto 0)) is
   begin
      
      out_trans.sig_CLK_out := signal_value;
      
   end procedure set_CLK;
   
   procedure set_CLK_oe          (signal_value : in std_logic) is
   begin
   
      out_trans.sig_CLK_oe := signal_value;
   
   end procedure set_CLK_oe;
   
   procedure get_DAT             (signal_value : out std_logic_vector(0 downto 0)) is
   begin

      signal_value := sig_DAT_in;
   
   end procedure get_DAT;
   
   procedure set_DAT             (signal_value : in std_logic_vector(0 downto 0)) is
   begin
      
      out_trans.sig_DAT_out := signal_value;
      
   end procedure set_DAT;
   
   procedure set_DAT_oe          (signal_value : in std_logic) is
   begin
   
      out_trans.sig_DAT_oe := signal_value;
   
   end procedure set_DAT_oe;
   
   procedure event_CLK_change is
   begin

      wait until (sig_CLK_in'event and out_trans.sig_CLK_oe = '0');

   end event_CLK_change;
   procedure event_DAT_change is
   begin

      wait until (sig_DAT_in'event and out_trans.sig_DAT_oe = '0');

   end event_DAT_change;

end altera_conduit_bfm_vhdl_pkg;

